Swedish translation of monotone - sv.po

The translation sv.po is distributed under the same license as
the monotone package.

Richard Levitte <richard@levitte.org>, 2006
Joel Rosdahl <joel@rosdahl.net>, 2006

Translation guidelines:
-----------------------
access                          åtkomst
address                         adress
ancestor                        förfader [eller förälder i vissa fall]
ancestry                        föräldraskap
approval                        godkännande
approve                         godkänna
argument                        argument
authenticate                    autentisera
author                          upphovsman
authorize                       auktorisera
automation                      automatisering
backup                          säkerhetskopia
bad                             felaktig
base (revision)                 grund(revision)
(to) bisect                     (att) dela upp
bisection                       uppdelning
bogus                           felaktig
bookkeeping directory           administrativ katalog
boolean                         boolesk
(a) branch                      gren
(to) branch                     förgrena
buffer                          buffert
bug                             fel / programfel
byte(s)                         byte()
cert(s)                         cert()
(a) change                      ändring
changelog (message)             loggmeddelande
(a) check                       kontroll
check out                       hämta
checksum                        kontrollsumma
child                           barn
client                          klient
(a) commit                      ändringar
(to) commit (to)                arkivera (i)
connect                         ansluta
connection                      anslutning
database schema                 databasschema
debug                           felsöka
default (foo)                   standard(foo)
delta                           delta
deny                            neka
descendent                      ättling
destination                     mål
directory                       katalog
disapproval                     underkännande
disapprove                      underkänna
disconnect                      koppla ifrån
divergence                      divergens
drop                            slänga / ta bort / överge
dump                            dumpa
edge                            båge
editor                          textredigerare
epoch                           epok
exchange                        utbyte
file                            fil
find                            leta
found                           hittade / hittat
get                             hämta
graph                           graf
(a) hash (value)                kontrollsumma
hash check                      kontrollsummering
head                            löv
history                         historik
host                            värd
hostname                        värdnamn
initialize                      initiera
(an) input                      indata
interface                       gränssnitt
invalid                         ogiltig
keystore                        nyckellager
log                             logg
malformed                       otydbart
manifest                        manifest
marking                         markering
(a) match                       matchning
(to) match (a pattern)          matcha
(to) match (a non-pattern)      stämma (med/överens)
(to) not match (a non-pattern)  skilja sig (ifrån) / inte stämma (med/överens)
(a) merge                       ihopslagning
(to) merge                      slå ihop
(log) message                   loggmeddelande
migrate                         migrera
migration                       migrering
(to) mismatch                   inte matcha / inte stämma överens
mismatched                      inkonsistent
node                            nod
(to) note                       notera
note:                           obs:
option                          flagga (i programanrop)
option                          inställning (i inställningsfiler)
output                          utmatning, utdata
(to) output                     (att) mata ut
(an) overflow                   överflöde
(to) overflow                   flöda över
override                        åsidosätta
packet                          paket
parent                          förälder
parse                           tyda
parseable                       uttydbar
parsing                         uttydning
passphrase                      lösen
path                            sökväg [eller fil/katalog i vissa fall]
pattern                         mönster
peer                            [formulera om]
(to) process                    behandla
progress                        förlopp
propagate                       propagera
pull                            hämta
push                            skicka
query                           fråga
rebuild                         bygga om
refined                         raffinerad
refuse                          neka
reject                          neka
repository                      arkiv
request                         begäran
revision                        revision
root                            rot
roster / rosters                lista / listor
selection                       val
selector                        väljare
serve                           servera
server                          server
service                         tjänst
(to) set                        sätta
sink                            mottagare
socket                          sockel
source                          källa
(to) specify                    (att) ange
specified                       angivna
stale                           trasig
state                           tillstånd
suspend                         avstängd / avstänga
sync                            synkronisera
synchronize                     synkronisera
tag                             tagg
terminate                       avbryta
tree                            träd
(an) underflow                  underflöde
(to) underflow                  flöda under
usher                           usher
violate                         ej uppfylla
work set                        arbetsmängd
workspace                       arbetskopia (el. kanske arbetskatalog, ibland)

If that isn't enough, maybe having a look at the swedish part of the
Translation Project might help:  http://www.tp-sv.se/
